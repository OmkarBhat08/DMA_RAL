class dma_agent extends uvm_agent;

	dma_sequencer seqr;
	dma_driver drv;
	dma_monitor mon;

	`uvm_component_utils(dma_agent)

	function new(string name = "dma_agent", uvm_component parent = null);
		super.new(name, parent);
	endfunction

	function void build_phase(uvm_phase phase);
		super.build_phase(phase);
		if(get_is_active() == UVM_ACTIVE)
		begin
			seqr = dma_sequencer::type_id::create("seqr", this);
			drv = dma_driver::type_id::create("drv", this);
		end
		mon = dma_monitor::type_id::create("mon", this);
	endfunction : build_phase

	function void connect_phase(uvm_phase phase);
		super.connect_phase(phase);
		drv.seq_item_port.connect(seqr.seq_item_export);
	endfunction : connect_phase

endclass : dma_agent
