class dma_test extends uvm_test;

	dma_env env;

	`uvm_component_utils(dma_test)

	function new(string name = "dma_test", uvm_component parent = null);
		super.new(name, parent);
	endfunction : new

	function void  
endclass : dma_test
